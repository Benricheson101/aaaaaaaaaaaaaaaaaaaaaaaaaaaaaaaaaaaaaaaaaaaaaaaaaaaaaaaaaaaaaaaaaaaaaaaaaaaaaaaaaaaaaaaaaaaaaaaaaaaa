module aaa(); 

initial begin
	forever begin
		$write("a")
	end
end

endmodule
